`include "mux2_1.v"

module mux2_1_tb;

    reg [31:0] in1, in2;
    reg s;

    wire [31:0] out;

    mux2_1 uut(in1, in2, s, out);

    initial
        begin
            $dumpfile("mux2_1_tb.vcd");
            $dumpvars(1, mux2_1_tb);
            
            #1
            s = 0;

            #1
            in1 = 32'b0000_0010_0000_0000_1111_0000_0000_1111;
            in2 = 32'b0010_0000_1111_0000_0000_0010_0000_0000;

            #1
            $display("out: %d", out);

            #1
            s = 1;

            #1
            in1 = 32'b0000_0010_0000_0000_1111_0000_0000_1111;
            in2 = 32'b0010_0000_1111_0000_0000_0010_0000_0000;

            #1
            $display("out: %d", out);

            #1
            s = 0;

            #1
            in1 = 32'b0010_0000_1111_0000_0000_0010_0000_0000;
            in2 = 32'b0000_0010_0000_0000_1111_0000_0000_1111;

            #1
            $display("out: %d", out);

            #1
            s = 1;

            #1
            in1 = 32'b0010_0000_1111_0000_0000_0010_0000_0000;
            in2 = 32'b0000_0010_0000_0000_1111_0000_0000_1111;

            #1
            $display("out: %d", out);

        end

endmodule