module image;

    reg [7:0] imfile [0:783]; // 28 * 28

endmodule