module instructionmemory(pc, instruction);

    input [9:0] pc; // change later
    
    output reg [31:0] instruction;

    reg [31:0] memfile [0:1023]; // increase memory size later

    initial
        begin // write instructions here
            // x0 = 0 already done

            //  addi x10, x0,  1
            //                immediate         rs1   func3   rd       opcode     
            memfile[0] <= 32'b0000_0000_0001___00000___000___01010___001_0011;          //  x10     =   1

            //  addi x11, x10, 1
            memfile[1] <= 32'b0000_0000_0001___01010___000___01011___001_0011;          //  x11     =   2

            //  addi x12, x10, 2
            memfile[2] <= 32'b0000_0000_0010___01010___000___01100___001_0011;          //  x12     =   3
              
            //  addi x13, x10, 3 
            memfile[3] <= 32'b0000_0000_0011___01010___000___01101___001_0011;          //  x13     =   4

            //  add  x14, x11, x13                                                                                               
            memfile[4] <= 32'b0000000___01011___01101___000___01110___011_0011;         //  x14     =   6   (x14 = x11 + x13)

            //  addi x15, x14, 0
            memfile[6] <= 32'b0000_0000_0000___01110___000___01111___001_0011;          //  x15     =   6   (x15 = x14 + 0)

            //  sub x16, x11, x15
            memfile[7] <= 32'b0100000___01011___01111___000___10000___011_0011;          // x16     =   4   (x16 = x15 - x11)

            //  addi x17, x16, 0
            memfile[8] <= 32'b0000_0000_0000___10000___000___10001___001_0011;          //  x17     =   4   (x17 = x16 + 0)

            //  sw   x11, 4(x0)         
            memfile[9] <= 32'b0000000___01011___00000___000___00100___010_0011;         //  mem[4]  =   2

            //  sw   x12, 5(x0)         
            memfile[10] <= 32'b0000000___01100___00000___000___00101___010_0011;         // mem[5]  =   3

            //  lw   x18, 5(x0)         
            memfile[11] <= 32'b0000_0000_0101___00000___000___10010___000_0011;         //  x18     =   mem[5] 

            //  addi x19, x18, 0
            memfile[12] <= 32'b0000_0000_0000___10010___000___10011___001_0011;          //  x19     =   3   (x19 = x18 + 0)

            //  addi x4, x3, 1
            //memfile[5] <= 32'b0000000___00000___00101___000___00101___000_0011;
        end

    always @ (pc)
        begin
            instruction <= memfile[pc];
        end

endmodule