module image;

    reg [45*7:0] imfile;

endmodule