module instructionmemory(pc, instruction);

    input [9:0] pc; // change later
    
    output wire [31:0] instruction;

    reg [7:0] memfile [0:1023]; // increase memory size later

    assign instruction = {memfile[pc+3], memfile[pc+2], memfile[pc+1], memfile[pc]};

    initial
        begin // write instructions here
            //  addi x10, x0,  1
            {memfile[3], memfile[2], memfile[1], memfile[0]} <= 32'b0000_0000_0000___00000___000___00000___001_0011;          //  x10     =   1

            //  addi x11, x10, 1
            {memfile[7], memfile[6], memfile[5], memfile[4]} <= 32'b0000_0000_0001___01010___000___00000___001_0011;          //  x11     =   2

            //  addi x12, x10, 2
            {memfile[11], memfile[10], memfile[9], memfile[8]} <= 32'b0000_0000_0010___01010___000___00000___001_0011;         //  x12     =   3

            //  nop
            {memfile[15], memfile[14], memfile[13], memfile[12]} <= 32'b0000_0000_0000___00000___000___00000___000_0000;        //  nop

            //  sw   x10, 9(x0)
            {memfile[19], memfile[18], memfile[17], memfile[16]}  <= 32'b0000000___01010___00000___010___01001___010_0011;       //  mem[9]  =   1

            //  nop
            {memfile[23], memfile[22], memfile[21], memfile[20]} <= 32'b0000_0000_0000___00000___000___00000___000_0000;        //  nop

            //  addi x13, x10, 3
            {memfile[27], memfile[26], memfile[25], memfile[24]} <= 32'b0000_0000_0011___01010___000___00000___001_0011;         //  x13     =   4

            //  add  x14, x13, x11 (rd, rs1, rs2)
            {memfile[31], memfile[30], memfile[29], memfile[28]} <= 32'b0000000___01011___01101___000___00000___011_0011;        //  x14     =   6   (x14 = x11 + x13)

            //  addi x15, x14, 0
            {memfile[35], memfile[34], memfile[33], memfile[32]} <= 32'b0000_0000_0000___01110___000___00000___001_0011;        //  x15     =   6   (x15 = x14 + 0)

            //  sub x16, x15, x11
            {memfile[39], memfile[38], memfile[37], memfile[36]} <= 32'b0100000___01011___01111___000___00000___011_0011;        // x16     =   4   (x16 = x15 - x11)

            //  addi x17, x16, 0
            {memfile[43], memfile[42], memfile[41], memfile[40]} <= 32'b0000_0000_0000___10000___000___00000___001_0011;        //  x17     =   4   (x17 = x16 + 0)

            //  sw   x11, 4(x0)
            {memfile[47], memfile[46], memfile[45], memfile[44]} <= 32'b0000000___01011___00000___010___00100___010_0011;       //  mem[4]  =   2

            //  nop
            {memfile[51], memfile[50], memfile[49], memfile[48]} <= 32'b0000_0000_0000___00000___000___00000___000_0000;       //  nop

            //  sw   x12, 5(x0)
            {memfile[55], memfile[54], memfile[53], memfile[52]} <= 32'b0000000___01100___00000___010___00101___010_0011;       // mem[5]  =   3

            //  nop
            {memfile[59], memfile[58], memfile[57], memfile[56]} <= 32'b0000_0000_0000___00000___000___00000___000_0000;       //  nop

            //  lw   x18, 5(x0)
            {memfile[63], memfile[62], memfile[61], memfile[60]} <= 32'b0000_0000_0101___00000___010___00000___000_0011;       //  x18     =   mem[5]  =   3

            //  nop
            {memfile[67], memfile[66], memfile[65], memfile[64]} <= 32'b0000_0000_0000___00000___000___00000___000_0000;       //  nop

            //  addi x19, x18, 0
            {memfile[71], memfile[70], memfile[69], memfile[68]} <= 32'b0000_0000_0000___10010___000___00000___001_0011;       //  x19     =   3   (x19 = x18 + 0)

            //  and  x20, x10, x18
            {memfile[75], memfile[74], memfile[73], memfile[72]} <= 32'b0000000___01010___10010___111___00000___011_0011;      //  x20     =   1   (x20 = x10 & x18)
            //  x10 = 0000_0000_0000_0000_0000_0000_0000_0001
            //  x18 = 0000_0000_0000_0000_0000_0000_0000_0011
            //  x20 = 0000_0000_0000_0000_0000_0000_0000_0001

            //  addi x23, x20, 0
            {memfile[79], memfile[78], memfile[77], memfile[76]} <= 32'b0000_0000_0000___10100___000___10111___001_0011;          //  x23     =   1   (x23 = x20 + 0)

            ///////////////////////
            //  or  x21, x11, x16
            {memfile[83], memfile[82], memfile[81], memfile[80]} <= 32'b0000000___01011___01111___000___00000___011_0011;       //  x21     =   6   (x21 = x11 | x16)
            //  x11 = 0000_0000_0000_0000_0000_0000_0000_0010
            //  x16 = 0000_0000_0000_0000_0000_0000_0000_0100
            //  x21 = 0000_0000_0000_0000_0000_0000_0000_0110

            //  addi x24, x21, 0
            {memfile[87], memfile[86], memfile[85], memfile[84]} <= 32'b0000_0000_0000___10101___000___00000___001_0011;       //  x24     =   6   (x24 = x21 + 0)

            //  xor  x22, x14, x17
            {memfile[91], memfile[90], memfile[89], memfile[88]} <= 32'b0000000___01110___10001___100___00000___011_0011;      //  x22     =   2   (x22 = x14 xor x17)
            //  x14 = 0000_0000_0000_0000_0000_0000_0000_0110
            //  x17 = 0000_0000_0000_0000_0000_0000_0000_0100
            //  x22 = 0000_0000_0000_0000_0000_0000_0000_0010

            //  addi x25, x22, 0
            {memfile[95], memfile[94], memfile[93], memfile[92]} <= 32'b0000_0000_0000___10110___000___00000___001_0011;      //  x25     =   2   (x25 = x22 + 0)

            //  nop
            {memfile[99], memfile[98], memfile[97], memfile[96]} <= 32'b0000_0000_0000___00000___000___00000___000_0000;      //  nop

            //  lw   x26, 4(x0)
            {memfile[103], memfile[102], memfile[101], memfile[100]} <= 32'b0000_0000_0100___00000___010___00000___000_0011;     //  x26     =   mem[4]  = 2

            //  addi x27, x26, 0
            {memfile[107], memfile[106], memfile[105], memfile[104]} <= 32'b0000_0000_0000___11010___000___00000___001_0011;      //  x27     =   2   (x27 = x26 + 0)

            //  nop
            {memfile[111], memfile[110], memfile[109], memfile[108]} <= 32'b0000_0000_0000___00000___000___00000___000_0000;      //  nop

            //  lw   x30, 9(x0)
            {memfile[115], memfile[114], memfile[113], memfile[112]} <= 32'b0000_0000_1001___00000___010___00000___000_0011;     //  x30     =   mem[9]  =   1

            //  nop
            {memfile[119], memfile[118], memfile[117], memfile[116]} <= 32'b0000_0000_0000___00000___000___00000___000_0000;     //  nop

            //  addi x31, x30, 0
            {memfile[123], memfile[122], memfile[121], memfile[120]} <= 32'b0000_0000_0000___11110___000___00000___001_0011;     //  x31     =   1

            //  sw   x24, 8(x16)
            {memfile[127], memfile[126], memfile[125], memfile[124]} <= 32'b0000000___11000___10000___010___00000___010_0011;   // mem[12]  =   6

            //  sw   x25, 9(x17)
            {memfile[131], memfile[130], memfile[129], memfile[128]} <= 32'b0000000___11001___10001___010___00000___010_0011;   // mem[13]  =   2

            //  sw   x19, 13(x10)
            {memfile[135], memfile[134], memfile[133], memfile[132]} <= 32'b0000000___10011___01010___010___00000___010_0011;   // mem[14]  =   3

            //  sw   x30, 12(x18)
            {memfile[139], memfile[138], memfile[137], memfile[136]} <= 32'b0000000___11110___10010___010___00000___010_0011;   // mem[15]  =   1

            //  lw   x5, 10(x11)
            {memfile[143], memfile[142], memfile[141], memfile[140]} <= 32'b0000000___01010___01011___010___00000___000_0011;   // x5   =   mem[12]  =   6

            //  lw   x6, 10(x12)
            {memfile[147], memfile[146], memfile[145], memfile[144]} <= 32'b0000000___01010___01100___010___00000___000_0011;   // x6   =   mem[13]  =   2

            //  lw   x7, 8(x15)
            {memfile[151], memfile[150], memfile[149], memfile[148]} <= 32'b0000000___01000___01111___010___00000___000_0011;   // x7   =   mem[14]  =   3

            //  lw   x8, 13(x25)
            {memfile[155], memfile[154], memfile[153], memfile[152]} <= 32'b0000000___01101___11001___010___01000___000_0011;        // x8   =   mem[15]  =   1

            //  addi x4, x5, 0
            {memfile[159], memfile[158], memfile[157], memfile[156]} <= 32'b0000_0000_0000___00101___000___00100___001_0011;         //  x5     =   6
            
            //  addi x4, x6, 0
            {memfile[163], memfile[162], memfile[161], memfile[160]} <= 32'b0000_0000_0000___00110___000___00100___001_0011;         //  x6     =   2

            //  addi x4, x7, 0
            {memfile[167], memfile[166], memfile[165], memfile[164]} <= 32'b0000_0000_0000___00111___000___00100___001_0011;         //  x7     =   3

            //  addi x4, x8, 0
            {memfile[171], memfile[170], memfile[169], memfile[168]} <= 32'b0000_0000_0000___01000___000___00100___001_0011;         //  x8     =   1
        end

endmodule