module convolution();

    reg signed [63:0] filter [0:2][0:2];

endmodule