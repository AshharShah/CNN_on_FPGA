module convolution();

    reg signed [31:0] filter [0:2][0:2];

endmodule