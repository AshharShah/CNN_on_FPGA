module image;

    reg [7:0] imfile [0:784];

endmodule