module image;

    reg [7:0] imfile [0:27][0:27]; // 28 * 28

endmodule