`include "alu.v"

module alu_tb;

reg [3:0] aluctl;
reg [31:0] a, b;
wire [31:0] out;
wire zero;
wire overflow;

alu          uutC(aluctl, a, b, out, zero, overflow);

initial
    begin
        $dumpfile("alu_tb.vcd");
        $dumpvars(1, alu_tb);

        // Testing AND function
        #1
        a       =   32'b0000_1111_0010_0000_0000_0110_0000_0011;
        b       =   32'b0000_1110_0010_0100_0100_0010_0000_0001;
        aluctl  =   4'b0000; // 0 AND

        #1
        $display("out 1: %d", out);

        #1
        a       =   32'b0000_1111_0000_1111_0000_1111_0000_1111;
        b       =   32'b1111_0000_1111_0000_1111_0000_1111_0000;
        aluctl  =   4'b0000; // 0 AND

        #1
        $display("out 1: %d", out);

        #1
        a       =   32'b1000_0000_1111_0000_0100_0000_0010_0001;
        b       =   32'b1000_0000_1111_0000_0010_0100_0010_0001;
        aluctl  =   4'b0000; // 0 AND

        #1
        $display("out 1: %d", out);

        //Testing OR function
        #1
        a       =   32'b1010_0000_1111_0010_0101_0010_0010_0001;
        b       =   32'b1010_0000_1111_1000_0011_0110_0010_0001;
                    //  1010_0000_1111_1010_0111_0110_0010_0001
        aluctl  =   4'b0001; // 1 OR

        #1
        $display("out 1: %d", out);

        #1
        a       =   32'b0000_0000_0000_0010_0111_0000_0010_0100;
        b       =   32'b0010_0010_1101_1010_0011_0111_0000_1001;
                    //  0010_0010_1101_1010_0111_0111_0010_1101
        aluctl  =   4'b0001; // 1 OR

        #1
        $display("out 1: %d", out);

        //Testing OR function
        #1
        a       =   32'b1010_0000_1111_0010_0101_0010_0010_0001;
        b       =   32'b1010_0000_1111_1000_0011_0110_0010_0001;
        //
        aluctl  =   4'b0010; // 2 ADD

        #1
        $display("out 1: %d + %d = %d", a, b, out);

        #1
        a       =   32'b0000_0000_0000_0010_0111_0000_0010_0100;
        b       =   32'b0010_0010_1101_1010_0011_0111_0000_1001;
        aluctl  =   4'b0010; // 2 ADD

        #1
        $display("out 1: %d + %d = %d", a, b, out);

        #1
        a       =   32'b1000_0000_1111_0000_0100_0000_0010_0001;
        b       =   32'b1000_0000_1111_0000_0010_0100_0010_0001;
        aluctl  =   4'b0010; // 2 ADD

        #1
        $display("out 1: %d + %d = %d", a, b, out);

        //Testing SUB function
        #1
        a       =   32'b1010_0000_1111_0010_0101_0010_0010_0001;
        b       =   32'b1010_0000_1111_1000_0011_0110_0010_0001;
        aluctl  =   4'b0110; // 6 SUB

        #1
        $display("out 1: %d - %d = %d", a, b, out);

        #1
        a       =   32'b0000_0000_0000_0010_0111_0000_0010_0100;
        b       =   32'b0010_0010_1101_1010_0011_0111_0000_1001;
        aluctl  =   4'b0110; // 6 SUB

        #1
        $display("out 1: %d - %d = %d", a, b, out);

        #1
        a       =   32'b1000_0000_1111_0000_0100_0000_0010_0001;
        b       =   32'b1000_0000_1111_0000_0010_0100_0010_0001;
        aluctl  =   4'b0110; // 3 SUB

        #1
        $display("out 1: %d - %d = %d", a, b, out);

        //Testing EQL function
        #1
        a       =   32'b1010_0000_1111_0010_0101_0010_0010_0001;
        b       =   32'b1010_0000_1111_1000_0011_0110_0010_0001;
        aluctl  =   4'b0111; // 7 EQL

        #1
        $display("out 1: %d == %d = %d", a, b, out);

        #1
        a       =   32'b0000_0000_0000_0010_0111_0000_0010_0100;
        b       =   32'b0010_0010_1101_1010_0011_0111_0000_1001;
        aluctl  =   4'b0111; // 7 EQL

        #1
        $display("out 1: %d == %d = %d", a, b, out);

        #1
        a       =   32'b1000_0000_1111_0000_0100_0000_0010_0001;
        b       =   32'b1000_0000_1111_0000_0100_0000_0010_0001;
        aluctl  =   4'b0111; // 7 EQL

        #1
        $display("out 1: %d == %d = %d", a, b, out);

        //Testing NOR function
        #1
        a       =   32'b1010_0000_1111_0010_0101_0010_0010_0001;
        b       =   32'b1010_0000_1111_1000_0011_0110_0010_0001;
        aluctl  =   4'b1100; // 12 NOR

        #1
        $display("out 1: %d", out);

        #1
        a       =   32'b0000_0000_0000_0010_0111_0000_0010_0100;
        b       =   32'b0010_0010_1101_1010_0011_0111_0000_1001;
        aluctl  =   4'b1100; // 12 NOR

        #1
        $display("out 1: %d", out);

        #1
        a       =   32'b1000_0000_1111_0000_0100_0000_0010_0001;
        b       =   32'b1000_0000_1111_0000_0100_0000_0010_0001;
        aluctl  =   4'b1100; // 12 NOR

        #1
        $display("out 1: %d", out);
    end

endmodule